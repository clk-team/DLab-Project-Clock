

module shower(
    input num,
    output a[7:0]
);