module musicwake(
   input do,
   output reg music
);