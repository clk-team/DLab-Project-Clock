`timescale 1ns/1ps

module set_time (
    
);

endmodule //set_time