module mode_selection(clk,sel);

input clk;
input [2:0]sel;

always@(posedge clk) begin
    

endmodule